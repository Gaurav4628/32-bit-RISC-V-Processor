`timescale 1ns / 100ps

module alu_ctrl(
    input [1:0] ALUOp,
    input [6:0] funct7,
    input [2:0] funct3,
    output reg [3:0] alu_ctrl
    );
    
    always@(*) begin
        case(ALUOp)
            2'b00 : alu_ctrl = 4'b0010; //load, store
            2'b01 : alu_ctrl = 4'b0110; // for branches
            2'b10 : begin
                case(funct3)
                    3'b000: begin
                        if(funct7 == 7'b0100000) alu_ctrl = 4'b0110; //SUB
                        else alu_ctrl = 4'b0010;
                        end
                    3'b111: alu_ctrl = 4'b0000; //AND
                    3'b110: alu_ctrl = 4'b0001; //OR
                    3'b010: alu_ctrl = 4'b0011; //SLT
                    3'b100: alu_ctrl = 4'b0010; //XOR 
                   default: alu_ctrl = 4'b0010;
                endcase
                end
             default: alu_ctrl = 4'b0010;
         endcase
         end
                 
endmodule

